/**
  @brief Memory Controller module that does memory controller controlling

  @note Interface is on nyu-ambam, which will be included as a package
*/
module MemCtrl(
  MemCommon_if.memCtrl mem 
);
  // Add memory controller logic here

endmodule
